��/      }��	Resultats�}�(�schema�]�(�Id��INT����Moyenne��FLOAT����Promo��INT����Grp��INT����Rang��INT���e�header_page_id�N�allocated_pages�]�(�managers.page_id��PageId���)��}�(�FileIdx�K �PageIdx�K ubh)��}�(hK hKubh)��}�(hK hKubh)��}�(hK hKubh)��}�(hK hKubh)��}�(hK hKubeus.